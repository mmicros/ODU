LIBRARY ieee;
USE ieee.std_logic_1164.all;
entity counter8 is
		port(x1: in std_logic;
			  f0, f1, f2, f3, f4, f5, f6, f7	 : out std_logic);
end counter8 ;

architecture count of slider is
signal cnt := 0;

begin 
	
end count;